`timescale 1ns / 1ps
module multiplexor(
    input  logic [3:0] user_input,   // usuario ingresa exactamente 4 bits
    output logic [6:0] display_out  // salida para display de 7 segmentos
);

    always_comb begin
     case (user_input)
     4'b0000: display_out = 7'b0000001;//#0
     4'b0001: display_out = 7'b1001111;//#1
     4'b0010: display_out = 7'b0010010;//#2
     4'b0011: display_out = 7'b0000110;//#3
     4'b0100: display_out = 7'b1001100;//#4
     4'b0101: display_out = 7'b0100100;//#5
     4'b0110: display_out = 7'b0100000;//#6
     4'b0111: display_out = 7'b0001111;//#7
     4'b1000: display_out = 7'b0000000;//#8
     4'b1001: display_out = 7'b0001100;//#9
     default: begin 
     display_out = 7'b1111111; // todo apagado si algo raro ocurre
     $display("Entrada inv�lida: %b", user_input);
     end           
     endcase
     end
     endmodule
